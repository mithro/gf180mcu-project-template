// SPDX-FileCopyrightText: © 2025 XXX Authors
// SPDX-License-Identifier: Apache-2.0

`default_nettype none

module chip_core #(
    parameter NUM_INPUT_PADS,
    parameter NUM_BIDIR_PADS,
    parameter NUM_ANALOG_PADS
    )(
    `ifdef USE_POWER_PINS
    inout  wire VDD,
    inout  wire VSS,
    `endif
    
    input  wire clk,       // clock
    input  wire rst_n,     // reset (active low)

    `ifndef MAX_IO_CONFIG
    input  wire [NUM_INPUT_PADS-1:0] input_in,   // Input value
    output wire [NUM_INPUT_PADS-1:0] input_pu,   // Pull-up
    output wire [NUM_INPUT_PADS-1:0] input_pd,   // Pull-down
    `endif

    input  wire [NUM_BIDIR_PADS-1:0] bidir_in,   // Input value
    output wire [NUM_BIDIR_PADS-1:0] bidir_out,  // Output value
    output wire [NUM_BIDIR_PADS-1:0] bidir_oe,   // Output enable
    output wire [NUM_BIDIR_PADS-1:0] bidir_cs,   // Input type (0=CMOS Buffer, 1=Schmitt Trigger)
    output wire [NUM_BIDIR_PADS-1:0] bidir_sl,   // Slew rate (0=fast, 1=slow)
    output wire [NUM_BIDIR_PADS-1:0] bidir_ie,   // Input enable
    output wire [NUM_BIDIR_PADS-1:0] bidir_pu,   // Pull-up
    output wire [NUM_BIDIR_PADS-1:0] bidir_pd   // Pull-down

    `ifndef MAX_IO_CONFIG
    ,inout  wire [NUM_ANALOG_PADS-1:0] analog  // Analog
    `endif
);

    // See here for usage: https://gf180mcu-pdk.readthedocs.io/en/latest/IPs/IO/gf180mcu_fd_io/digital.html

    `ifndef MAX_IO_CONFIG
    // Disable pull-up and pull-down for input
    assign input_pu = '0;
    assign input_pd = '0;
    `endif

    // Set the bidir as output
    assign bidir_oe = '1;
    assign bidir_cs = '0;
    assign bidir_sl = '0;
    assign bidir_ie = ~bidir_oe;
    assign bidir_pu = '0;
    assign bidir_pd = '0;
    
    logic _unused;
    assign _unused = &bidir_in;

    logic [NUM_BIDIR_PADS-1:0] count;

    // Count increments when all input bits are set (or always if no inputs)
    wire count_enable;
    `ifdef MAX_IO_CONFIG
    assign count_enable = 1'b1;  // Always count when no inputs (MAX_IO_CONFIG)
    `else
    generate
        if (NUM_INPUT_PADS > 0) begin : gen_count_enable
            assign count_enable = &input_in;
        end else begin : gen_count_enable_default
            assign count_enable = 1'b1;  // Always count when no inputs
        end
    endgenerate
    `endif

    always_ff @(posedge clk) begin
        if (!rst_n) begin
            count <= '0;
        end else begin
            if (count_enable) begin
                count <= count + 1;
            end
        end
    end

    logic [7:0] sram_out;

    gf180mcu_fd_ip_sram__sram512x8m8wm1 sram (
        `ifdef USE_POWER_PINS
        .VDD  (VDD),
        .VSS  (VSS),
        `endif

        .CLK  (clk),
        .CEN  (1'b1),
        .GWEN (1'b0),
        .WEN  (8'b0),
        .A    ('0),
        .D    ('0),
        .Q    (sram_out)
    );

    assign bidir_out = count ^ {{(NUM_BIDIR_PADS-8){1'b0}}, sram_out};

endmodule

`default_nettype wire
